---------------------------------------------------------------------------------
-- This is free and unencumbered software released into the public domain.
--
-- Anyone is free to copy, modify, publish, use, compile, sell, or
-- distribute this software, either in source code form or as a compiled
-- binary, for any purpose, commercial or non-commercial, and by any
-- means.
--
-- In jurisdictions that recognize copyright laws, the author or authors
-- of this software dedicate any and all copyright interest in the
-- software to the public domain. We make this dedication for the benefit
-- of the public at large and to the detriment of our heirs and
-- successors. We intend this dedication to be an overt act of
-- relinquishment in perpetuity of all present and future rights to this
-- software under copyright law.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
-- EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE AUTHORS BE LIABLE FOR ANY CLAIM, DAMAGES OR
-- OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
-- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
-- OTHER DEALINGS IN THE SOFTWARE.
--
-- For more information, please refer to <http://unlicense.org/>
---------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity rom_40x128_exclif1_ip is
    port (
        clka : in std_logic;
        addra : in std_logic_vector(5 downto 0);
        douta : out std_logic_vector(767 downto 0)
    );
end entity rom_40x128_exclif1_ip;

architecture behavior of rom_40x128_exclif1_ip is


    type rom_type is array (0 to 40) of std_logic_vector(767 downto 0);


    constant mem : rom_type := (
"000011000011000010000011000000000101000000111101111101111110000001000010111101000000000011111110111110000000000000111101111101000000111101111110000001000010111110000001000001111111000100000010111101111100111110000101000011000011000000000001000000000001000001111011000001111111000000000001000110000000111101000010111111111110000010000000111110111100111101000001111111000000111111111111000000000011111101111110000001000011000001000110000000000001111100000001000010000000000010111111000001111111000011111110000001000011000001111011000011111110111101000010000000000011111111111110000101111100111101111100000000000000111011000011000000000011111111000000000011000000000000000000111110111110111110111101111011111111000000111110000000000010000000000001000000000001111111111101",
"111110111111000101000000000000111111000000000000111011111101111110111100000000000001000010111101000011111111000010111101111101000001000010111101000010111101111111000001111111000100111110111101000001111111000010000001111100000000111011111111000101000011111110111100111010000100111110111110000000111110111101000100000100000011000100111110000010111101000000111010000100000011000000111100111101111100000000000001111110000010000101111110000001000000111110111111000010111111000010000010111110111100111011000011000000111110000011000000111101111101111110111111000100000000111111111101000010000000000000000100000100000000000001111110000011000001000000000101000011000000000100000011111101000100000000000001000100111111111111000100000011111111000010111011000100111101111101000011",
"000001111111000101000001000100111110000000000000111011111111000100111100111111000011000000111110111110111110111110111010000001000000000100000011111101000010000000000011000011000101111110000011000010000000111100000011000001111101111100000010111111111111111100000010111110000101111111000000111110000011000101111101111010111110000100000010000010000000000100111111111111111011111100111111000010111100111110111101000000000010000010000001000010111111111111000011000001000100111100000100000010111101111110000100000001000100000101111111000010111101111110000000000010000100111111000000111110000011111111111111111111000000111100111010000000111101111111000000111111000011111101000100111100000001000000000010000100000011111101000011000011111110111101111101111100111111000000000000",
"111111111111000000000001111110111101111111111100000001000000000010000011000101000010000010000100000000111101000110111101000010000100111111000000000000000000000010000010000100000001000100111101000011111101000010000000000000000000111110111010000010000010000001111101111101000100111110111101000011111101000101000010111010000010000010000011111101000100000010110111111100000001000011111101000101000001111111000000000001000000000000111110000100111110000000000001000000000100000000000101111101111111110111000100000001111110111111000100000000111110111100000000000101000100000010000000111110000000000000000000111111000011000000111100000011000011000010000000111110000000000100111110111101111111111111000000000000111110000010111111000001000000000011111110000000111011000011111110",
"000011000011000000111111111100000101000100111100000010000011000011000011000100000000000011000000000011000011000000111010000101000011111100000001111111000010111101111110111100000001000000000100111100111101111111111100000001111010111101111001111101000010111111111101111110111110000000111111111101000101000000111101111101000000000000111111111110111011000000111000000000111011000000000000000000111010000000000000111101000000000011000101000101000000000100000001000001000000000000111111000000111011111001000001000000111111000010000010111111111001000010000000111110000100000110000010111110111111000011000001000010000001000001000011000011000101000100000001111101000011000001111101111111000001111111111101111011000100000000000000000011111111111101000010000000000010000000000100",
"111111000010111111000100000100000001000000000000000000111011000001000011000011000000000100000010000011000010111111111100000000000011000000000001000010000010000000111111000000000000000011000000111111000001111110000100111100000010111101111110000100000001111001111110111100111111000001000100111110000000111111111111111101111111000101000011000011111101000101111001111111000010111110000001111101111110111100000000000000000001111101000101000000111110000100000100000011111101000100111110000001111101111000000010111101000000000011111110000001000001111111000100111101000001000000000001000101000001000001000010111110000000000001111111000011000001000000000001000000000100000101000000000000111110111011000000000000111111111111000000000011000001000011111101000000111110000100111111",
"000001000001111011000011000011111111000001000100111111000000000101000000000010111101000001000011000000000100111110111010111110000000000000000000000000111111111110000100111101111110000110111101000001000011111010111101111111000010000010111110000000000000111100111101111010000001000000000001111111000010111111000000111110000101000010111010000000000011000001111100000001000011000000000001111111000000111111000001000010000011000011111101111011000000000100000011000101111110000011000001000100111101111011000001000110000000111110111111000000111111111100000011111100000000000010000011000010000010111100111111000101000010000000111100111011000101000011111111111110000001000001000001000010000011000000000100000000111110000100000000000011000011000000000100000001000011000000000100",
"000001000010000001000000000100000011000100111110000101111110000000000011000001110111111011000101111110000000000110111010000101111101000100111110111111000001000100111101111101111111111111000101000010000011000000000000111110000000000010111011000100000000111111111100111111000101111100111111001000000010111100000010111011000011000101111000000011000100000110111010000010111101111010000011000000000100111110111111000010111111111010111110111001111100111101000010000011000001000001000010000010000001111110000011000011000011111101000011111111111111000010000000000011111111111110000000000110000011111110111010000000111111000011111110000000000001000000111010000001111100111101111011111110111110000001111110000101111110111100111001111010000101000000000000111100111100000101000110",
"000100000011000011000100111110111100000011000001111111000100000000000000111011111110111101000101000000111111001000111111000000111111000101000001111111111100000011000000111110000000111110000010000110111111111011000011000000111011000010111101000000111111000001000011111011000000111101000010000010000111000001000100111111000001111111111010000100111110111110111001000000000000111101111101111101000101000001111100111011111110111100111101111010111010000000000000111110001000000110000010111110111111111101000010000101000111111011000011000000000000000011111111000000000000000101000101000000000100000010111110111111111101000101111001000000111100111011000000000000000000111100111001111111111101111111111011000011111100111100111011000001000010111011000100000001000000111101000000",
"000010000001111101111111000000111101111111000101000010111101000000000010111111110111000000000101000000110111000000111101000011111110000101111100111010000000000000000000000000000111000100000011000110111111000001000000000000000011111110111110111110111111111110000010000001111011000011000101000101000110000010000101111110000101000011111001000001000000000000000011000001000011111010111110000000000000000000111010111111000000000000111101000010111011111111000001000110000100000000000001000000000010111110111111000101000011111101000000111110000011111101000000000000111100000000000011000100000101111111111101111110111010000001000000000101111011111111000000000000111101000001000000111110000001000011000000000011111100111010111001111010000110000001000000111011111100000010000000",
"111110111100000000000000000011000001000011000011000101111110000010000110000100111010111101000001111111111010000011000001000010000010000001000001111110000010000011111111111111000011000110000101000010000011000011000000000001000000111101000000111111000100000001000011111011111011111010000010000101000000000100111101111111111101000100111001000011000001000000111011000000000010111111111100000001000001111011000000000010111010111011000000000001111111000001000100000010111111000101000010001000111100000011000110000001111111111101000000000001111100000100000110000011111101111000000100000000111110111111000000000100000011000000000100000000000000111110000010000010000001111011000010111111000001111101000000000000000101111011111001111110000111111010000001111101000000000000000000",
"000000000000000000000000111100000000000100000011111110000001000101000000000110000000000010111100111111111010000001111101111111111011000011111011111011111111111110000000000001111101111100111110111100111100111011111011111111111101111101000000000001111111111100111110111110111101000000000000111110111101000100000000111110111111111110000000111100000000000100111001111011000000000001000011000001000010000001000011000000000000111111000100111011111111111010111110000000111011000001111110000111000000000110000110111110000000111100111101111011111110000000111110111101111101111010000001000001111111000000111100000101111110000000000010111101111010111111111110111010111100000001111100000010111111000000000001000100000111111110111110111111111110111011000101000011000000000110000010",
"000000111111000001111101111110000001000011000000000101000010000011000000111111000000000011000001000100000000000100000000000010111110000001000000111111111111000110000001111111111010111110000000000010000000000000000010111110000011111111000101000000111111111101000010111110000111000000000011111101111100000001000100111101000000000011000010000100000011000110111010000000000011000010000001000000000100000001111110111111000101000001000011111110000011000000000001000101111010000110000000000000000000000000111110000100111001111111000101000100000001111110111100111101000010111011000000000000000001111011000011000001000101000101000010111010000011000000000010111110000000111101000001000011111100000001111111000000000111000101000100111101111101000001000010000000000101000010111001",
"111110111111000010111110000100000001111110000000000011111110000010111101000100000011111101111101111100000100000001000001111111111111111100000011111111000000000001111110000011111110111001111111000110000001111011111111111100111111000000111100000100111101111111000000111011000101000100111011111110111101000001111100000011111100111110111110111011111111000000000000111101000011000100000000000011000000111010000010000001000100000010000001111111000010111111000010111101111101000011111111000100111100111101000100000010111110000011000000111111000000111101111110111010111110111101111100000100000110000001111101111101111111000110000100111110111100000100000000111011000001111110111100000001000010111101000000111100000011000110000001111111111101000001000000000000111111000010111010",
"000000000000111100000000111111111111000101000010000000000010111100111101000101000011000010000000000011000011111110111110111110000000111101000010000010111110111111000100000001111010111110000000111101000100000001000001111010111011111110111101111111000000111010000010000000000000000001111100000100111111111101000011000000000000111011111111000000000100111100000001111101111110000010000101111110111110000000000101000011111110111111000001000000000101000100000001111101000000000001000000000101111111000001111100000001000001111100111100111111111011111111000010000000000101111111111101111011000000111000000010111100000110000000000101111111111111000011000101000100111101000011000001111101000101000000111100111100000010000000000011111100000100000010111011000000111011000100111110",
"000011000100111111000100000101000110111111111111111100000010111101111101111111000000000001111111111011000100111100111110111111000010000001000000000010111111111110111111111111111111111100000001111100000011111011000011111110111111000100111000111101000001110111000000111001000100000011000010000000111111111110000001000000111100111100111001000000000101000011111110000000000011000011000010000000000001000001000101000000000101000011000100000000000101000011000010000001111111111011111110000000000011111000111110111110000001111101111111000110000000000101111111111100000110111101111101000010000010000000111110000000000100111110000101111111000001000101000100000000111011000011000000111101111111111110111100000010000010000010000010111100111101000000111101000000111110111100111110",
"111101111110111100111101000010000001000001111110111110111011111100000000000011000100000010111100111100000000111111111110000000000010000000000001000100000010111111000110111110111101111110111101111101000001000010000000000010000010111110111001000010111100111001000100000001000110000001000110000000111011000000000010000001111100000100111001111111000010111101111011111100000001000100000101000110000010111100000000000000111111111110000110000010000101000000111110000000111100111111111101000010000010111001111011000010000001000010000101000110111100000011000001111101000010000100000000000000000001111101000001000011111110111111000000111110000100000101111100000011111111111110000101111110111110000000000100000010111110000101000000111101111011111111000000111100111010111101000011",
"000011111110000000000101111111000011111100000011000110000000111011111100000010000000111100000011000000000000000010111101111111000000000110000000000000000011000110000110111100111010111110000001000011000010000000000001111000111110111100111011000000000000111111000011000010000001000001000010000110111011000001111101111111111111111111111011000100111110111101000010111100111111000010111111000010000000111111000010111111000011111101000000111100111110000001000011111010000001000000000010111101111111000000000000000000111011000100000011000001111111000000111111000000000000000000000100111111000001000000111111000100111111111101111110111100000101111101111101111111111101000010000011000001000000000000111011000100000001000000000111000010111101000000000000000001111100111110000000",
"000001000000111101111110000100000000111100000010000011111110111101111110111110000010000000000010111111000011111101111111111110111101111111111110000010111101000000000001000011000000000011111101111111111111000100000010111011111110111110111101000001000010000001000100111011000001000000000111000110000000000111000101111110000001111000111011111100000001111010111111000000000001000000111111000011000100000001111110111110111101000000000001000010111111000000111110111010111100111101000010111100000000111111111110111111000000111110000010000010111011000100000000111000000001000000111111111100111100111010000011000000000011000010000011111101000101000010000010000011000001000001000100111101000011111011000011000100111100000010000000111101000001111111000000111100111011111101000011",
"000011000100000001111110000011000000111111111011111110111011111111000011111111000000000000111110000000000000000011111110000001111110000001000000000101000000111110000010111011111100000001000010000000000000000100000100111010111010000000111101000000111111000000000011000011000000000010000000000001000010000100000000111111000100111011111100111001000000000011000001000000000101000110000011000001000100111110000110000000111101111101111101000010000011000100000000111100000010000010111011111100111101000001111111111101000001111111000000000101111100000000000101111100000000000011000100000000000001111001000001111011000000000011000011000010000000000000000000000011111111000001000000000100000000111101000011000011000001000110000111000100111101000101000001000011111001000010111100",
"000000111111111111111111111111000010111011111110000011111111111111000011000000000101000001000010000001000000111110000100000010000001000011000011111111111111000000000000000001000001000000000010111110111100000000000101000010000011000001111101000100000000111011000011111110000100000011111101000000111100000110000001111111111110111110000100000000000101111101000100111111111101111111111111111101000010000010000000000000000000111111000011000001000100000000111111111111000000000010111110111001000000000000111101000000111011000100111110000100000000000101111100111110000010000011000010000000000000111100000001111100000101000100111111000011000011111111000100000001111111000101000000000000000011000000000000000000111101111111111111111101000000000000000001111111000010111101000000",
"000001111100111110111111000110111110111100000100000100111110000011111010111111000010000011000001111101111111000010000100111110000000111101000110000000000010000011000001111101111111000001000001000000111100000100000110111101111101111111000001000000111100111111000010000011000011111111000000111110000000000110111011000000111011111101000000111110000000111110000000000011111110000100000011000100000001111101000010000100000010000010111111000011000001000100000001111100111100111011000100000001111011000000000001000000000000000011000000000111000000000010111011111110000011000000000001000000111101111111000011000000000100000100111111111110000110111110000001000100000010000011000010000100000001000000000000000100000000000010111111000011111100000010111100000011111101111011111100",
"000011111100111100000000111111000000111110000011000011000000111111000001111101000011000100111100000100000000111100111101000000111101111110111111000010000101000000111101000100111101111100000011000011000100111101000010000000111100000001000000111010000000111111000001000000000100000010000001000001000010000101111100000001111000000000000100000101111111000101000000000100000001000011000001111010000000111110111110111111000000111100000110000001000011111101111110111101111100000010111100111110111111000001111101000101111101111100111111000000000111000000000011111110000110111111000011111001111101111111111110000011111011111111111111111110000000000010000011000011111110000100000101000000000111000000000100111100111100000000000000000001111000000100111111000100000101111011000000",
"111100111010000000000001000011111110111111000010000001111101000011111101000110000011000010111011000001000111111100000011000100000010111110000011000000000000000011111011000101000100000011000101000101000010000010000000000101000101000000000010111100000001111101111111000101111110000000000000111101000000111011111001111111111001000011000101000010111111000000000100000011000011000110111110111010000001000000111111000001000100111111000001000010000000111110111111111110111110000000000100111110111011000101000000000001000000111110111111000101000000000000111110000011000100000010111100111100111010000011000011000010111011000001000000111110001000000101000010000000000100000001000100000001000100000001000101000000111010000000000001111111000000000001000000000011000101111010111110",
"000010000000111011111110000110111001111110000110000110111110000000111100000000111110000001111111000010000001000010000001000100000000111010000010000011000100111111111101000110111101000001000000000101000010000000111011000110000001111011000111000000000011000101000000000001000000111111111010111110111111111011111010111111111001111111000010000101000000000000000100000111111111000000000101111100000011000000000110000010000100000001000110000011111101000010000001000001000000111100000000111100000011000010000000000110000001111101000011000000000010111101111111000001000100001000000001111000000010000000000000111010111110000101111110000000000101111101000011000011000101000010000111111110000110000101111111111100000011111111000001000011000011001000000001111100000000111000111110",
"111110000000111100000000111110111011111110111101111111111101000010000000000011000110111100111001000110000000111111000000111110000101111001111110000010000000000000000000000010111110111110000111000010000011000010111111000011111110000000000000000001111111000000000010000010000000000011111010111001111100111101000000000001110111000001000001001000111011111101000101000000111100111110000110111010000010000000000011000011000010000000000011000001111110000000111010000101111011111011111110111100111100000001000011000100111111111001000100111111000000000001000110000110001000000100000001111001000001000000111111111101111100000001000011000010000001000100111111000010000101111111000000000100000001111111000101111111000000000000000101111101000001000110000000000000000101111011000100",
"000000111101000000111001000010111010000001000010000001111111111111111001111111000011000001000000000001001000111100000000000000111110111001000010111101111101000001111100000100000100111101000010000110111101111111111001000010111110000010000111111100111101000000000000000101111010000100111111111001111011000010111100000000111011111011000111000011000001111110000000000101111101000100000100000001000000111110000000000001000011111011000111111111111110111111111100000011111101000001000000111001111100000100000001000001000110111101000011000101000101000010111111000000000101000110000000111000000000000111000011000001111111000011000000111100000001000000000010000001000001111101000000000011111111111111000000111001111110000010000011000010000000000110000000000100111110111000111111",
"111111111100111111111011000100111100111101000000000000111011000011111011000000000000111111111011000011111111000010000010111111000000111101000101000010111100000001111100000000000010000100000110000011000000000011111011111110000010000010000000000001000000000010000001000100111111111100111011111100000010000000111100000010111101111111000000000110111101000010111101000000000011000110000010111010111111000000000101000100111101111010000011000001111111111100111100111110000010111111111110111011111110000001000000000111000000000001111101000111000110000001000000000010000110000000111111111101111110000101000011111111111110000101000001111011111101000001000011111100000010111111000110000101111110000101000000111100111010000101000110111111000010000111000010000001000000111110000100",
"000011111011111111111111000000111010111011000000000110111110111111111001000000000011000000000001000001000101000010000000000110000100111111000011000011000010111101111011000000111110111101000001000110111101111111111010000001000000111101111111111001111111000000000010000001111100000000111110111010000100111100111001000000000000111110111111111111111110111111000101000010111100000000000000111010000000000010111111000010111011000001000100111111000011111101111100111110000100111100000010000000111110000000000010000001000010111101000100000011000111000011000100111110000010000010000000111101111101000101111111000000000001000001111110111110000101000000111110111011000001000000000001000010111100000000000001111011111010111101000001111111000000000110111100000000000010111001000000",
"000000111101111110111011000101000010111100111111000000111110000011000000111110000000000010111010000000000100000010000000000101111110000001000011111110000011111111111101111111000000111111000000000010000001000000000001111111000101000010000000111010000010000101000000000000000000000000000101000000000001000011111100000011000000111110000010000000000001111100000000000100000000000010000110000101000010000011000011000010000000111111000000000001000001000000111101000000000101111101000101000000111100000101111101000011000101111110111101000000000000111101000110000101000011000001111110000001111100000010000010111101111011111110000010000000000010000010000010111111000011000000000111111111111110000010000001111011000000111101111110111011000110111111111101000000000111111010000011",
"000000000010111110111010000100111011111010000000000011111011000000000010111100000011111110111101000100000001111100000011111111111101111110000000000010000000000000000010000101000010000100111110000110000010000000111101000100111110000000000100111010000010000110000100111110111110000001000111000011000000000010000000000010000001000011000010001000111110111100000001111111000001111101111111000000000000111010000011111110111111111101000000111111000101000011000000000010000101111111000010111111000010000000000000000111000000111011000000000000111111111110000000000011000001000010111101000000111001000101000010000001111010000010000100111110000001111011111111111100000010000000000111000000111111000110000001000000000100111111000010111111111110000110000001000100000000111001000100",
"111101000010000011111110000101111110111111000110000100000010111011111111000010000000111101111000000101000000000000000100111110000000000000111110000000111110000000000011000000111101000001000000000101111110000000111111000001000101111111001000111101000000000000111101000000000010000000000100000101111111111111111010111110111111000011000001000010000001000010000000000000000010000011000100000111000000111100000100000000111100000001000011000011111111000000111011111110111101000000000000000010000001000110111100000000000110111110111100000101000000000100000000000000000100000000111011000100111110000000000000111100111100000000000001000010111110000000111101000010111011111111000001000101111010111111000001111111000100000100000000111111111110000011000011111111000011000001111111",
"000000000010000001111100000101111111111000000100000010111110111011111101111011000101000000111010111111000100000001000000000011000001111011000011000010111011000001000010111101000010111111000100000101000110000100000000000011000001000000000000111111111110000010111111000100111010111101000000000000000100000010111011000000000010111110000001000111111011000000000101000011000101000001000100000110000101111110000011000011111011111101000001000000000001000001000001000011111111000110000001111110000001000011111011000010000111111101000100000010111101000011000001000000000000111101000000000011111110000010111101111101111100000101000010000000000100111111111111111100111110000100111110000101111011000101111110111101000011000010000001111010000101000000000100000000000110111111000011",
"111100111111000000111010000000000001111010000100000110111101111011000000111100000000111101000001111100000100000000000000000101000100000000000001111110111010000010000001000011111110000100000110000000111111000011000001111110000101000011000000111011111101000100000001111101111100000100000001000001111110111100111110111100000001000100000000000101000010000000000100111111111110000000111111000011000010000000000011111111111100111101000110000000000011000000111101000000000100000101111111000000111100000101111111111111111111111110111101000110111100000000000001111011000000111101111100000001111101111111111101111111111011111111000011111011111101000000111101111110000001000000111101000000111111000100000000111111000000111110000101000010000000000010000101111111000011000100000000",
"111110000000000100111011000010111010000000111111000001000000111110000101000010111111000101111011111101111111000000111101000100111100111111000000000000111111001000000010000000111100000000111101000101000000000000000000000000111110000001000011111110111011111110000000000010000001000000000100000001000010000000111101000100111101000100000000000010000011111111000001000000000000000001111101111111000100111011000010111111111101000011000011000000000011000000000011000011000100000001000000000000111011000001111111000010000000111111000010000110111111111110001000000000000000111111111100000100000000000100000010111100111101000110000000000000111111111110000001000000111111000000000001111100000000000011000010111101111111000110111111111010000000000001000100111111111110000110000000",
"000000000100000001111001000000000000111010000010000010111110111111000001000001000011000010111001000011111101000000000000000010000100111110000011111101111011111111000101111101111011000110000011000010111110000011000001000010111111111101000101111110111011000011111111111101111100000001000010000001000001000000111111111101000000000101000010000000000101000100111110000011000000000011000010000110111111111100000010111100111110111111000011000000111110000010111101000000111111000100111101111111000001000001111111000010000110111110111101000100111110111110000001111110000000111111000000000011000000000100111010000000111100000000000001111110000011111011111110000000000000000001111111111101000000111111111111000100000001111110000000111001000001000000000000111110111111000010000010",
"000100000000000110000010000011111101111100111101000101111111111111000100111110000001111110111111111111000011000100000101000110111101000001111111111101111011000011000001000000000000000000000011000000000000000001000001000011000100111111111111000000000000000100000001000001000001000000000011000000000101111100111100111110000000000101111101000110000001000001000011111101111110000100111111000000000000000010000100000100000000111100000000000000000110111111000001000000000101000010111111111110111111111110000001000011000010111101000000000000111011000001000011111110111101000000000010000000000011111100111110111101111001000101000010111101000001000010000000000000000000000010111011000000111100111111000001000011000100000011000100000000000011111111000000000011111110111111000011",
"000011111110000010111101000000111011000001000000000000000011000000000101000010000000000000111001111100000010111111000000000000111111111100000010000000111011000001000011000010000010000011111110000100000011000011000000111110111100111110000100000000111110111111000000111101000011111111000000000100000000000000000101000001000001000001000100000000000011111110111100111101000001000011111101000100000001000000000001000000000010000001000001000100000001000000111110000100111110000100000000000010000000000010111011111111111111111100111101000001111100000001000111000000111110111010111010000101000100000000000000000010111001111111111111111101111100111010111111111101000001111111111110000010000000000011000100000101000101000011000000000000000000111100000001111111000000000100000101",
"111111000010000100000010111110111101111101000000000010111101111100111110111101000001000000000000000001111110111110000101000011111110000011000011000100000010111110000100000011000100000101111111000101000000000001000001111011000011000000000110000010000001000011000000000001111100000000000010000101000000000000111110000001000000000100000011000001000001000000000000111101111101111111111110000001000001111111000000111110000000111110111101111111111101000000000011000100000010111101111111000010000100000000000000000000000101111111000010111110111010000000000000000011111011111111000001000100000011111111000011000000000011000011111101000101111100111101000010000010000001000000000001000100111011000001000000000101111101000011000101000001000010111111111111111100000000000100000100",
"000000000000111111000010000011000011000100111110000011000001000101111101000100000100000010111100000000000001111101000100000010000000000000000000000100111111111100000100000010000000111110000100000000000001000011000000000000000100000000111100000000000100000000111101111100111011000000000010111111000000000000000000111111000000111111111111111101111101000000111111111111000000000011111100000010111110111111000011111101000011000000111110000011000010111111111110111111000001111101111111000001000001000010000000111110000000111101000000111101000000111110000000000100000101111111000001000001111110000010000100111110000010111110000010111110111101000000111110000000111100000100000001000010000011000000111101111100000100111110000011111101000011111100000001000001000000000100111100",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");

begin

    rom_behavior : process(clka )
    begin

        if clka'event and clka='1' 
        then

            douta <= mem(to_integer(unsigned(addra)));

        end if;

    end process rom_behavior;


end architecture behavior;

