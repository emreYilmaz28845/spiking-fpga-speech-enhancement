---------------------------------------------------------------------------------
-- This is free and unencumbered software released into the public domain.
--
-- Anyone is free to copy, modify, publish, use, compile, sell, or
-- distribute this software, either in source code form or as a compiled
-- binary, for any purpose, commercial or non-commercial, and by any
-- means.
--
-- In jurisdictions that recognize copyright laws, the author or authors
-- of this software dedicate any and all copyright interest in the
-- software to the public domain. We make this dedication for the benefit
-- of the public at large and to the detriment of our heirs and
-- successors. We intend this dedication to be an overt act of
-- relinquishment in perpetuity of all present and future rights to this
-- software under copyright law.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
-- EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE AUTHORS BE LIABLE FOR ANY CLAIM, DAMAGES OR
-- OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
-- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
-- OTHER DEALINGS IN THE SOFTWARE.
--
-- For more information, please refer to <http://unlicense.org/>
---------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity rom_128x10_exclif2_ip is
    port (
        clka : in std_logic;
        addra : in std_logic_vector(6 downto 0);
        douta : out std_logic_vector(59 downto 0)
    );
end entity rom_128x10_exclif2_ip;

architecture behavior of rom_128x10_exclif2_ip is


    type rom_type is array (0 to 128) of std_logic_vector(59 downto 0);


    constant mem : rom_type := (
"111101000010111111000000000000000010111101111111000000000011",
"000011000000111011111111000011000000000001111100111101000000",
"111010111100000010000001000000000010000010111100111010000010",
"111101000000000000000000000000000010111111000001111111000010",
"000000000000000000000000000100000000000000000000111111000000",
"111100000011000000000001111101000000111111000000111011000010",
"111110111100111111000000111111000011000011111110111110000011",
"111111111111000000111111111101111110000000111111000000000000",
"111011000000111101000001111110111101000011000001111000000100",
"111110000000111111000000000000111110000011000101111100000000",
"000001111100000000111111000001000000000100000000111111000010",
"000000000001111110111110000001000000111111111110000000000000",
"111110111111111111000000111110000000111111000000000000000000",
"111101111111000100000010000001000000000001111100111101000000",
"000010000010111111000000111111111100111110111011111110000010",
"111100111011000011000000111111000010000000000000111101111101",
"111100000011000001000001111101111100000011000000000000000010",
"000000000000111111000000111111111111000001000010111110000000",
"111110111110000001111111111101111101000001000010000000000001",
"000000000001111111111111000000000001111111111111111111000001",
"000011000000111111000000111011111011111111000010000001000000",
"000000000000111111000000000000111101111111000000000000000011",
"111111000011000000000001111111111101000001111111000000111111",
"000000000000111111000000111111000001111111000000000010000000",
"111000111011000000111111000000000110000100000100110111111111",
"000010111110000011000000000000111111111101000001111111111101",
"000011000000111111000000111110111100000011111111000000000001",
"111111111110000000111110000011000000000010000000000010000001",
"111111111111111111000000000000111110000000000000000000000010",
"111011111111000001000000111101000000111110111001111000000010",
"000010111111000000111100000010000000000000111110111110000000",
"000010111101111111111110000001000010111111000000000001111110",
"000001000001111110111111000000111110111100111110000011000000",
"111001000011000000111111110111000000111111111100111011000000",
"000000000010000001000010111111111101000000000000000000000000",
"000000111111000001000001111100000001111011000000000001000110",
"111100111111111101111111111111000010000000000001111100000000",
"000000111101000000111101000001000000111100000011111110111111",
"111010111101000011000000111101111110111110111010111100111111",
"111110000001111110000010000000000000000000000010111110111110",
"111111000000000010111101000000000000000000111101000000111110",
"000100111111111111111110111101111111000011000000000001111101",
"111101000000000000000001000000000101000001000000000000000000",
"000000000000000010000001111111000010111101000000111110111111",
"000010111101000010111100111111111111111110000010000011000001",
"111011110111000010000000000010000010000001111101110110111111",
"000000000000000000111110111111000000000001000000000010000001",
"000000111011111110111011000000111111000010111110000000000011",
"000001111110000010000000111110000000000000000000000000111111",
"000001111101000001000000000011000001000001000000000010000000",
"111100111111111110000000000000000011111110000000000001000001",
"000000111110000010000000000010000001000000000010000001000010",
"000001000000000000111111111111000001000000111110000000111111",
"111111000010111101000010000001000000000011111111111110000010",
"111110111111111011111111111101000000000010000100111010000000",
"000010000000111101111111111010111011000000000011111110000001",
"000000000000000010000010000000111101000010000000000000000000",
"000100111100000000111100000000111100000001000000000000111100",
"000001000001000001000001000000111111000000000000000001000010",
"111111000000000000000000111110000001000000000001000000000010",
"111101000000111111000001111110000001000001000011111110000000",
"000000000000111111111111111111111111111110000000000000111111",
"111111000000000010111101000001000000000000000001000000111011",
"111111000000111100111101000001000010000010111010111101111110",
"111100000000000001000010111110111101000001000010111101111111",
"000000000000000000000000111110111101000000000100111101000001",
"000000111111000000111111000000000001000011000001000010111111",
"111101000001000011000001111101000000000000111111111100000001",
"111100111100000100000000000010000000000001000001111011111111",
"111111111011000001111010000000111110111101000000000000000000",
"000010000010111111111110000001111110111110000001000000111111",
"111011000000000001000000000001000001000000000000111100000010",
"111011111100000010000010111101000000000000111111111001000110",
"000000111110000001000000000010000010111110000010111111000000",
"000000000000111010111011111111000010111110111110000001111110",
"111111000000000010111110111111111111000010000001000000000000",
"000000111111111101111110000000000001000001111101000010000000",
"000001000001000000000000000000111101000000000000000010111111",
"111110111101111110111100111101000001111100000000000000000000",
"000000000010111101111011000000000001111111111101000000111110",
"000000000000111011111010000001000101000001000000000001111110",
"111110000001000000000000000000111111000000000100111101000000",
"000000000000000001000000000000111101000000111101000000111111",
"111110111110000011000010000000000000000001000010111111000010",
"111111000001000001111110000001111111000000000100111111111111",
"111001111000000010111111000100111111000000111001111100000000",
"000000000000000001111101111111000000000000111110000000000011",
"000000111111111111111100111111111110000000111111000000111111",
"111010111000000010000000000011000000000100111000111011000010",
"000000000000111111000000000000000000000000000000111101000001",
"000000111110000010000000000000000011000100111101111111000000",
"111011111101000010000010000000111110000001111100000000000011",
"000000000010111110111110000000111111000000000000000000111111",
"111100111101000010111111000000000010111111000100111100000001",
"111110000000000000000000000000000000000010000000000000111110",
"000001000001000010000001000001000011000000000001111111111111",
"111110000000111111000000000000000001111110000000000000000000",
"111101000001000000111110000000000001000000000100000000000001",
"111111111001111101111101111010000000111111000001000010000011",
"000011000000000000000011111100111111000000111111111110000010",
"111111000000111110000000000000111101000000111111000000111101",
"000001111111000001111111000011000000000000111011000000111011",
"000000000000111110000001000000111101111111111101000001000001",
"111110000010111100000000111110000000000000000000111100000100",
"111101000000111111000001000000000000111110000010000000000000",
"000001000000111101111111000001000000111111111101000011000000",
"111111000000000000000000111110000000000010000000000000000000",
"111110000001000000000000000000000000111101000001000000000000",
"111111111110000101111110000001000010111110111011111110000000",
"000001111100000000111100000001000000111100000000000000111110",
"111010000000111111000001111111000001000000000011111000000010",
"000001000000000010000000111101000000000000111111111110000000",
"000010111110111101111110111110000000111100000000000011000000",
"000001000000000001000001000000000000000001000010000001000000",
"111100000000111110000000111111000000000010000000111010000011",
"000010111111000010111110000001111110000000000001111111000011",
"000000111100111011111111000010000010111111000001000010000010",
"000000111111000010111111000001111111111110000010000011000010",
"000001111110000000111110111111000000111110000000111110000000",
"111111111111000000000000000010111111111111111110111111111011",
"111100111111000011000000000010000001000000111111111110000000",
"000001111101111111111110000001000000000000111111000000000011",
"000000000010111111111101000000000000000011111111111111000000",
"111110000001111111000000000000000000000000000000111110000000",
"000001000000111111111111000001000000000000111111000000000001",
"000001111101000010111011111111000000000001000010000000111100",
"000010000001111101111100111111000010000000000010000001000000",
"111111000010000010111110111110000001000010111111000010000000",
"000000000000000000000000000000000000000000000000000000000000");

begin

    rom_behavior : process(clka )
    begin

        if clka'event and clka='1' 
        then

            douta <= mem(to_integer(unsigned(addra)));

        end if;

    end process rom_behavior;


end architecture behavior;

